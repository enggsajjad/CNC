;
-- note PWMGenOutA = PWM, PWMGenOutB = DIR, PWMGenOutC = ENA

QuadB(1) <= IOBits(0);
QuadA(1) <= IOBits(1);
QuadB(0) <= IOBits(2);
QuadA(0) <= IOBits(3);
Index(1) <= IOBits(4);
Index(0) <= IOBits(5);
AltData(6) <= PWMGenOutA(1);
AltData(7) <= PWMGenOutA(0);
AltData(8) <= PWMGenOutB(1);
AltData(9) <= PWMGenOutB(0);
AltData(10) <= PWMGenOutC(1);
AltData(11) <= PWMGenOutC(0);
QuadB(3) <= IOBits(12);
QuadA(3) <= IOBits(13);
QuadB(2) <= IOBits(14);
QuadA(2) <= IOBits(15);
Index(3) <= IOBits(16);
Index(2) <= IOBits(17);
AltData(18) <= PWMGenOutA(3);
AltData(19) <= PWMGenOutA(2);
AltData(20) <= PWMGenOutB(3);
AltData(21) <= PWMGenOutB(2);
AltData(22) <= PWMGenOutC(3);
AltData(23) <= PWMGenOutC(2);

QuadB(5) <= IOBits(24);
QuadA(5) <= IOBits(25);
QuadB(4) <= IOBits(26);
QuadA(4) <= IOBits(27);
Index(5) <= IOBits(28);
Index(4) <= IOBits(29);
AltData(30) <= PWMGenOutA(5);
AltData(31) <= PWMGenOutA(4);
AltData(32) <= PWMGenOutB(5);
AltData(33) <= PWMGenOutB(4);
AltData(34) <= PWMGenOutC(5);
AltData(35) <= PWMGenOutC(4);
QuadB(7) <= IOBits(36);
QuadA(7) <= IOBits(37);
QuadB(6) <= IOBits(38);
QuadA(6) <= IOBits(39);
Index(7) <= IOBits(40);
Index(6) <= IOBits(41);
AltData(42) <= PWMGenOutA(7);
AltData(43) <= PWMGenOutA(6);
AltData(44) <= PWMGenOutB(7);
AltData(45) <= PWMGenOutB(6);
AltData(46) <= PWMGenOutC(7);
AltData(47) <= PWMGenOutC(6);

QuadB(9) <= IOBits(48);
QuadA(9) <= IOBits(49);
QuadB(8) <= IOBits(50);
QuadA(8) <= IOBits(51);
Index(9) <= IOBits(52);
Index(8) <= IOBits(53);
AltData(54) <= PWMGenOutA(9);
AltData(55) <= PWMGenOutA(8);
AltData(56) <= PWMGenOutB(9);
AltData(57) <= PWMGenOutB(8);
AltData(58) <= PWMGenOutC(9);
AltData(59) <= PWMGenOutC(8);
QuadB(11) <= IOBits(60);
QuadA(11) <= IOBits(61);
QuadB(10) <= IOBits(62);
QuadA(10) <= IOBits(63);
Index(11) <= IOBits(64);
Index(10) <= IOBits(65);
IOBits(66) <= PWMGenOutA(11);
IOBits(67) <= PWMGenOutA(10);
IOBits(68) <= PWMGenOutB(11);
IOBits(69) <= PWMGenOutB(10);
IOBits(70) <= PWMGenOutC(11);
IOBits(71) <= PWMGenOutC(10);

QuadB(13) <= IOBits(72);
QuadA(13) <= IOBits(73);
QuadB(12) <= IOBits(74);
QuadA(12) <= IOBits(75);
Index(13) <= IOBits(76);
Index(12) <= IOBits(77);
IOBits(78) <= PWMGenOutA(13);
AltData(79) <= PWMGenOutA(12);
AltData(80) <= PWMGenOutB(13);
AltData(81) <= PWMGenOutB(12);
AltData(82) <= PWMGenOutC(13);
AltData(83) <= PWMGenOutC(12);
QuadB(15) <= IOBits(84) ;
QuadA(15) <= IOBits(85) ;
QuadB(14) <= IOBits(86);
QuadA(14) <= IOBits(87);
Index(15) <= IOBits(88);
Index(14) <= IOBits(89);
AltData(90) <= PWMGenOutA(15);
AltData(91) <= PWMGenOutA(14);
AltData(92) <= PWMGenOutB(15);
AltData(93) <= PWMGenOutB(14);
AltData(94) <= PWMGenOutC(15);
AltData(95) <= PWMGenOutC(14);
