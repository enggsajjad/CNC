module aa(q,c,g);
    input q;
    input c;
    output g;



endmodule
